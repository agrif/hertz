// The below text was generated automatically by hertz
// using the {skeleton_name} skeleton.

module {toplevel_entity}();

endmodule
